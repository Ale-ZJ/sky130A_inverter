** sch_path: /home/alexandra/inverter/xschem/inverter_tb.sch
**.subckt inverter_tb out in
*.opin out
*.opin in
x1 net1 out in GND inverter
V1 in GND PWL(0 0 20n 0.0 900n 1.8)
.save i(v1)
V2 net1 GND 1.8
.save i(v2)
**** begin user architecture code

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


.control
save all
tran 1n 1u
plot v(in) v(out)
.endc

**** end user architecture code
**.ends

* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/alexandra/inverter/xschem/inverter.sym
** sch_path: /home/alexandra/inverter/xschem/inverter.sch
.subckt inverter vdd out in vss
*.iopin vdd
*.iopin vss
*.opin out
*.ipin in
XM1 out in vss vss sky130_fd_pr__nfet_01v8 L=0.18 W=4.5 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.18 W=3 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
