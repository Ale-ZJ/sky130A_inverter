magic
tech sky130A
magscale 1 2
timestamp 1671837334
<< error_p >>
rect -29 181 29 187
rect -29 147 -17 181
rect -29 141 29 147
rect -125 -147 -67 -141
rect 67 -147 125 -141
rect -125 -181 -113 -147
rect 67 -181 79 -147
rect -125 -187 -67 -181
rect 67 -187 125 -181
<< nwell >>
rect -311 -319 311 319
<< pmos >>
rect -114 -100 -78 100
rect -18 -100 18 100
rect 78 -100 114 100
<< pdiff >>
rect -173 88 -114 100
rect -173 -88 -161 88
rect -127 -88 -114 88
rect -173 -100 -114 -88
rect -78 88 -18 100
rect -78 -88 -65 88
rect -31 -88 -18 88
rect -78 -100 -18 -88
rect 18 88 78 100
rect 18 -88 31 88
rect 65 -88 78 88
rect 18 -100 78 -88
rect 114 88 173 100
rect 114 -88 127 88
rect 161 -88 173 88
rect 114 -100 173 -88
<< pdiffc >>
rect -161 -88 -127 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 127 -88 161 88
<< nsubdiff >>
rect -275 249 -179 283
rect 179 249 275 283
rect -275 187 -241 249
rect 241 187 275 249
rect -275 -249 -241 -187
rect 241 -249 275 -187
rect -275 -283 -179 -249
rect 179 -283 275 -249
<< nsubdiffcont >>
rect -179 249 179 283
rect -275 -187 -241 187
rect 241 -187 275 187
rect -179 -283 179 -249
<< poly >>
rect -33 181 33 197
rect -33 147 -17 181
rect 17 147 33 181
rect -33 131 33 147
rect -114 100 -78 126
rect -18 100 18 131
rect 78 100 114 126
rect -114 -131 -78 -100
rect -18 -126 18 -100
rect 78 -131 114 -100
rect -129 -147 -63 -131
rect -129 -181 -113 -147
rect -79 -181 -63 -147
rect -129 -197 -63 -181
rect 63 -147 129 -131
rect 63 -181 79 -147
rect 113 -181 129 -147
rect 63 -197 129 -181
<< polycont >>
rect -17 147 17 181
rect -113 -181 -79 -147
rect 79 -181 113 -147
<< locali >>
rect -275 187 -241 283
rect 241 187 275 283
rect -33 147 -17 181
rect 17 147 33 181
rect -161 88 -127 104
rect -161 -104 -127 -88
rect -65 88 -31 104
rect -65 -104 -31 -88
rect 31 88 65 104
rect 31 -104 65 -88
rect 127 88 161 104
rect 127 -104 161 -88
rect -129 -181 -113 -147
rect -79 -181 -63 -147
rect 63 -181 79 -147
rect 113 -181 129 -147
rect -275 -249 -241 -187
rect 241 -249 275 -187
rect -275 -283 -179 -249
rect 179 -283 275 -249
<< viali >>
rect -241 249 -179 283
rect -179 249 179 283
rect 179 249 241 283
rect -17 147 17 181
rect -161 1 -127 71
rect -65 -71 -31 -1
rect 31 1 65 71
rect 127 -71 161 -1
rect -113 -181 -79 -147
rect 79 -181 113 -147
<< metal1 >>
rect -253 283 253 289
rect -253 249 -241 283
rect 241 249 253 283
rect -253 243 253 249
rect -29 181 29 187
rect -29 147 -17 181
rect 17 147 29 181
rect -29 141 29 147
rect -167 71 -121 83
rect -167 1 -161 71
rect -127 1 -121 71
rect 25 71 71 83
rect -167 -11 -121 1
rect -71 -1 -25 11
rect -71 -71 -65 -1
rect -31 -71 -25 -1
rect 25 1 31 71
rect 65 1 71 71
rect 25 -11 71 1
rect 121 -1 167 11
rect -71 -83 -25 -71
rect 121 -71 127 -1
rect 161 -71 167 -1
rect 121 -83 167 -71
rect -125 -147 -67 -141
rect -125 -181 -113 -147
rect -79 -181 -67 -147
rect -125 -187 -67 -181
rect 67 -147 125 -141
rect 67 -181 79 -147
rect 113 -181 125 -147
rect 67 -187 125 -181
<< properties >>
string FIXED_BBOX -258 -266 258 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 0.18 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc +40 viadrn -40 viagate 100 viagb 0 viagr 0 viagl 0 viagt 100
<< end >>
